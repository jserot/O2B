custom-gcd.vhd