ENTITY __entity_name IS PORT(
  signal clk : IN STD_LOGIC; -- CPU's master-input clk (required for multi-cycle)
  signal reset : IN STD_LOGIC; -- CPU's master asynchronous reset (required for multi-cycle)
  signal clk_en: IN STD_LOGIC; -- Clock-qualifier (required for multi-cycle)
  signal start: IN STD_LOGIC; -- True when this instr. issues (required for multi-cycle)
  signal done: OUT STD_LOGIC; -- True when instr. completes (required for variable muli-cycle)
  signal dataa: IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- operand A (always required)
  signal datab: IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- operand B (optional)
  signal n: IN STD_LOGIC_VECTOR (7 DOWNTO 0); -- N-field selector (required for extended)
  signal a: IN STD_LOGIC_VECTOR (4 DOWNTO 0); -- operand A selector (used for Internal register file access)
  signal b: IN STD_LOGIC_VECTOR (4 DOWNTO 0); -- operand B selector (used for Internal register file access)
  signal c: IN STD_LOGIC; -- result destination selector (used for Internal register file access)
  signal readra: IN STD_LOGIC; -- register file index (used for Internal register file access)
  signal readrb: IN STD_LOGIC; -- register file index (used for Internal register file access)
  signal writerc: IN STD_LOGIC; -- register file index (used for Internal register file access)
  signal result : OUT STD_LOGIC_VECTOR (31 downto 0) -- result (always required)
END __entity_name;
