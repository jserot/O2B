-- platform.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity platform is
	port (
		altpll_0_areset_conduit_export    : in    std_logic                     := '0';             --    altpll_0_areset_conduit.export
		altpll_0_locked_conduit_export    : out   std_logic;                                        --    altpll_0_locked_conduit.export
		button_external_connection_export : in    std_logic_vector(1 downto 0)  := (others => '0'); -- button_external_connection.export
		clk_clk                           : in    std_logic                     := '0';             --                        clk.clk
		hex0_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   hex0_external_connection.export
		hex1_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   hex1_external_connection.export
		hex2_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   hex2_external_connection.export
		hex3_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   hex3_external_connection.export
		hex4_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   hex4_external_connection.export
		hex5_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   hex5_external_connection.export
		led_external_connection_export    : out   std_logic_vector(9 downto 0);                     --    led_external_connection.export
		reset_reset_n                     : in    std_logic                     := '0';             --                      reset.reset_n
		sdram_clk_clk                     : out   std_logic;                                        --                  sdram_clk.clk
		sdram_wire_addr                   : out   std_logic_vector(12 downto 0);                    --                 sdram_wire.addr
		sdram_wire_ba                     : out   std_logic_vector(1 downto 0);                     --                           .ba
		sdram_wire_cas_n                  : out   std_logic;                                        --                           .cas_n
		sdram_wire_cke                    : out   std_logic;                                        --                           .cke
		sdram_wire_cs_n                   : out   std_logic;                                        --                           .cs_n
		sdram_wire_dq                     : inout std_logic_vector(15 downto 0) := (others => '0'); --                           .dq
		sdram_wire_dqm                    : out   std_logic_vector(1 downto 0);                     --                           .dqm
		sdram_wire_ras_n                  : out   std_logic;                                        --                           .ras_n
		sdram_wire_we_n                   : out   std_logic;                                        --                           .we_n
		switch_external_connection_export : in    std_logic_vector(9 downto 0)  := (others => '0')  -- switch_external_connection.export
	);
end entity platform;

architecture rtl of platform is
	component platform_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component platform_altpll_0;

	component platform_button is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component platform_button;

	component platform_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component platform_cpu;

	component platform_hex0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component platform_hex0;

	component platform_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component platform_jtag_uart;

	component platform_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component platform_led;

	component platform_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component platform_onchip_memory;

	component platform_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component platform_sdram;

	component platform_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component platform_switch;

	component platform_sys_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component platform_sys_timer;

	component platform_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			led_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                       : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                      : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                             : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                         : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                                : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			button_s1_address                                          : out std_logic_vector(1 downto 0);                     -- address
			button_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_address                                : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                  : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                   : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                            : out std_logic;                                        -- debugaccess
			hex0_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			hex0_s1_write                                              : out std_logic;                                        -- write
			hex0_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex0_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			hex0_s1_chipselect                                         : out std_logic;                                        -- chipselect
			hex1_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			hex1_s1_write                                              : out std_logic;                                        -- write
			hex1_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex1_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			hex1_s1_chipselect                                         : out std_logic;                                        -- chipselect
			hex2_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			hex2_s1_write                                              : out std_logic;                                        -- write
			hex2_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex2_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			hex2_s1_chipselect                                         : out std_logic;                                        -- chipselect
			hex3_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			hex3_s1_write                                              : out std_logic;                                        -- write
			hex3_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex3_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			hex3_s1_chipselect                                         : out std_logic;                                        -- chipselect
			hex4_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			hex4_s1_write                                              : out std_logic;                                        -- write
			hex4_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex4_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			hex4_s1_chipselect                                         : out std_logic;                                        -- chipselect
			hex5_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			hex5_s1_write                                              : out std_logic;                                        -- write
			hex5_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex5_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			hex5_s1_chipselect                                         : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                          : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                           : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                     : out std_logic;                                        -- chipselect
			led_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                               : out std_logic;                                        -- write
			led_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                                          : out std_logic;                                        -- chipselect
			onchip_memory_s1_address                                   : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory_s1_write                                     : out std_logic;                                        -- write
			onchip_memory_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect                                : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                                     : out std_logic;                                        -- clken
			sdram_s1_address                                           : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                             : out std_logic;                                        -- write
			sdram_s1_read                                              : out std_logic;                                        -- read
			sdram_s1_readdata                                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                         : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                        : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                     : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                       : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                        : out std_logic;                                        -- chipselect
			switch_s1_address                                          : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_timer_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			sys_timer_s1_write                                         : out std_logic;                                        -- write
			sys_timer_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_timer_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			sys_timer_s1_chipselect                                    : out std_logic                                         -- chipselect
		);
	end component platform_mm_interconnect_0;

	component platform_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component platform_irq_mapper;

	component platform_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component platform_rst_controller;

	component platform_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component platform_rst_controller_002;

	signal altpll_0_c0_clk                                               : std_logic;                     -- altpll_0:c0 -> [cpu:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:altpll_0_c0_clk, onchip_memory:clk, rst_controller_002:clk, sdram:clk, sys_timer:clk]
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(26 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(26 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest             : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                 : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                     : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                    : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                   : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                    : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                      : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                      : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_sys_timer_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	signal mm_interconnect_0_sys_timer_s1_readdata                       : std_logic_vector(15 downto 0); -- sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	signal mm_interconnect_0_sys_timer_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	signal mm_interconnect_0_sys_timer_s1_write                          : std_logic;                     -- mm_interconnect_0:sys_timer_s1_write -> mm_interconnect_0_sys_timer_s1_write:in
	signal mm_interconnect_0_sys_timer_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                           : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                        : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                               : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                      : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                              : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_led_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                             : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                                : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_button_s1_readdata                          : std_logic_vector(31 downto 0); -- button:readdata -> mm_interconnect_0:button_s1_readdata
	signal mm_interconnect_0_button_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_s1_address -> button:address
	signal mm_interconnect_0_switch_s1_readdata                          : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_hex0_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	signal mm_interconnect_0_hex0_s1_readdata                            : std_logic_vector(31 downto 0); -- hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	signal mm_interconnect_0_hex0_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex0_s1_address -> hex0:address
	signal mm_interconnect_0_hex0_s1_write                               : std_logic;                     -- mm_interconnect_0:hex0_s1_write -> mm_interconnect_0_hex0_s1_write:in
	signal mm_interconnect_0_hex0_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	signal mm_interconnect_0_hex1_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	signal mm_interconnect_0_hex1_s1_readdata                            : std_logic_vector(31 downto 0); -- hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	signal mm_interconnect_0_hex1_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex1_s1_address -> hex1:address
	signal mm_interconnect_0_hex1_s1_write                               : std_logic;                     -- mm_interconnect_0:hex1_s1_write -> mm_interconnect_0_hex1_s1_write:in
	signal mm_interconnect_0_hex1_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	signal mm_interconnect_0_hex2_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	signal mm_interconnect_0_hex2_s1_readdata                            : std_logic_vector(31 downto 0); -- hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	signal mm_interconnect_0_hex2_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex2_s1_address -> hex2:address
	signal mm_interconnect_0_hex2_s1_write                               : std_logic;                     -- mm_interconnect_0:hex2_s1_write -> mm_interconnect_0_hex2_s1_write:in
	signal mm_interconnect_0_hex2_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	signal mm_interconnect_0_hex3_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	signal mm_interconnect_0_hex3_s1_readdata                            : std_logic_vector(31 downto 0); -- hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	signal mm_interconnect_0_hex3_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex3_s1_address -> hex3:address
	signal mm_interconnect_0_hex3_s1_write                               : std_logic;                     -- mm_interconnect_0:hex3_s1_write -> mm_interconnect_0_hex3_s1_write:in
	signal mm_interconnect_0_hex3_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	signal mm_interconnect_0_hex4_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	signal mm_interconnect_0_hex4_s1_readdata                            : std_logic_vector(31 downto 0); -- hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	signal mm_interconnect_0_hex4_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex4_s1_address -> hex4:address
	signal mm_interconnect_0_hex4_s1_write                               : std_logic;                     -- mm_interconnect_0:hex4_s1_write -> mm_interconnect_0_hex4_s1_write:in
	signal mm_interconnect_0_hex4_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	signal mm_interconnect_0_hex5_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	signal mm_interconnect_0_hex5_s1_readdata                            : std_logic_vector(31 downto 0); -- hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	signal mm_interconnect_0_hex5_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex5_s1_address -> hex5:address
	signal mm_interconnect_0_hex5_s1_write                               : std_logic;                     -- mm_interconnect_0:hex5_s1_write -> mm_interconnect_0_hex5_s1_write:in
	signal mm_interconnect_0_hex5_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- sys_timer:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:led_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal cpu_debug_reset_request_reset                                 : std_logic;                     -- cpu:debug_reset_request -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_002_reset_out_reset_req                        : std_logic;                     -- rst_controller_002:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sys_timer_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_sys_timer_s1_write:inv -> sys_timer:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv               : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_led_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_hex0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex0_s1_write:inv -> hex0:write_n
	signal mm_interconnect_0_hex1_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex1_s1_write:inv -> hex1:write_n
	signal mm_interconnect_0_hex2_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex2_s1_write:inv -> hex2:write_n
	signal mm_interconnect_0_hex3_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex3_s1_write:inv -> hex3:write_n
	signal mm_interconnect_0_hex4_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex4_s1_write:inv -> hex4:write_n
	signal mm_interconnect_0_hex5_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex5_s1_write:inv -> hex5:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [button:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, led:reset_n, switch:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n, sdram:reset_n, sys_timer:reset_n]

begin

	altpll_0 : component platform_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                 -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => sdram_clk_clk,                                  --                    c1.clk
			areset             => altpll_0_areset_conduit_export,                 --        areset_conduit.export
			locked             => altpll_0_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c2                 => open,                                           --           (terminated)
			c3                 => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	button : component platform_button
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button_s1_address,          --                  s1.address
			readdata => mm_interconnect_0_button_s1_readdata,         --                    .readdata
			in_port  => button_external_connection_export             -- external_connection.export
		);

	cpu : component platform_cpu
		port map (
			clk                                 => altpll_0_c0_clk,                                   --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	hex0 : component platform_hex0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex0_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_hex0_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_hex0_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_hex0_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_hex0_s1_readdata,           --                    .readdata
			out_port   => hex0_external_connection_export               -- external_connection.export
		);

	hex1 : component platform_hex0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex1_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_hex1_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_hex1_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_hex1_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_hex1_s1_readdata,           --                    .readdata
			out_port   => hex1_external_connection_export               -- external_connection.export
		);

	hex2 : component platform_hex0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex2_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_hex2_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_hex2_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_hex2_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_hex2_s1_readdata,           --                    .readdata
			out_port   => hex2_external_connection_export               -- external_connection.export
		);

	hex3 : component platform_hex0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex3_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_hex3_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_hex3_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_hex3_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_hex3_s1_readdata,           --                    .readdata
			out_port   => hex3_external_connection_export               -- external_connection.export
		);

	hex4 : component platform_hex0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex4_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_hex4_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_hex4_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_hex4_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_hex4_s1_readdata,           --                    .readdata
			out_port   => hex4_external_connection_export               -- external_connection.export
		);

	hex5 : component platform_hex0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex5_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_hex5_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_hex5_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_hex5_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_hex5_s1_readdata,           --                    .readdata
			out_port   => hex5_external_connection_export               -- external_connection.export
		);

	jtag_uart : component platform_jtag_uart
		port map (
			clk            => altpll_0_c0_clk,                                               --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	led : component platform_led
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,             --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv,     --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,           --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,          --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,            --                    .readdata
			out_port   => led_external_connection_export                -- external_connection.export
		);

	onchip_memory : component platform_onchip_memory
		port map (
			clk        => altpll_0_c0_clk,                               --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_002_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_002_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	sdram : component platform_sdram
		port map (
			clk            => altpll_0_c0_clk,                                 --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	switch : component platform_switch
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,          --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,         --                    .readdata
			in_port  => switch_external_connection_export             -- external_connection.export
		);

	sys_timer : component platform_sys_timer
		port map (
			clk        => altpll_0_c0_clk,                                --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_sys_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                        --   irq.irq
		);

	mm_interconnect_0 : component platform_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                            => altpll_0_c0_clk,                                           --                                          altpll_0_c0.clk
			clk_clk_clk                                                => clk_clk,                                                   --                                              clk_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			cpu_reset_reset_bridge_in_reset_reset                      => rst_controller_002_reset_out_reset,                        --                      cpu_reset_reset_bridge_in_reset.reset
			led_reset_reset_bridge_in_reset_reset                      => rst_controller_001_reset_out_reset,                        --                      led_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                    => cpu_data_master_address,                                   --                                      cpu_data_master.address
			cpu_data_master_waitrequest                                => cpu_data_master_waitrequest,                               --                                                     .waitrequest
			cpu_data_master_byteenable                                 => cpu_data_master_byteenable,                                --                                                     .byteenable
			cpu_data_master_read                                       => cpu_data_master_read,                                      --                                                     .read
			cpu_data_master_readdata                                   => cpu_data_master_readdata,                                  --                                                     .readdata
			cpu_data_master_write                                      => cpu_data_master_write,                                     --                                                     .write
			cpu_data_master_writedata                                  => cpu_data_master_writedata,                                 --                                                     .writedata
			cpu_data_master_debugaccess                                => cpu_data_master_debugaccess,                               --                                                     .debugaccess
			cpu_instruction_master_address                             => cpu_instruction_master_address,                            --                               cpu_instruction_master.address
			cpu_instruction_master_waitrequest                         => cpu_instruction_master_waitrequest,                        --                                                     .waitrequest
			cpu_instruction_master_read                                => cpu_instruction_master_read,                               --                                                     .read
			cpu_instruction_master_readdata                            => cpu_instruction_master_readdata,                           --                                                     .readdata
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,              --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                 --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,             --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,            --                                                     .writedata
			button_s1_address                                          => mm_interconnect_0_button_s1_address,                       --                                            button_s1.address
			button_s1_readdata                                         => mm_interconnect_0_button_s1_readdata,                      --                                                     .readdata
			cpu_debug_mem_slave_address                                => mm_interconnect_0_cpu_debug_mem_slave_address,             --                                  cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                  => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                                     .write
			cpu_debug_mem_slave_read                                   => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                                     .read
			cpu_debug_mem_slave_readdata                               => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                                     .readdata
			cpu_debug_mem_slave_writedata                              => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                                     .writedata
			cpu_debug_mem_slave_byteenable                             => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                                     .byteenable
			cpu_debug_mem_slave_waitrequest                            => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                                     .waitrequest
			cpu_debug_mem_slave_debugaccess                            => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                                     .debugaccess
			hex0_s1_address                                            => mm_interconnect_0_hex0_s1_address,                         --                                              hex0_s1.address
			hex0_s1_write                                              => mm_interconnect_0_hex0_s1_write,                           --                                                     .write
			hex0_s1_readdata                                           => mm_interconnect_0_hex0_s1_readdata,                        --                                                     .readdata
			hex0_s1_writedata                                          => mm_interconnect_0_hex0_s1_writedata,                       --                                                     .writedata
			hex0_s1_chipselect                                         => mm_interconnect_0_hex0_s1_chipselect,                      --                                                     .chipselect
			hex1_s1_address                                            => mm_interconnect_0_hex1_s1_address,                         --                                              hex1_s1.address
			hex1_s1_write                                              => mm_interconnect_0_hex1_s1_write,                           --                                                     .write
			hex1_s1_readdata                                           => mm_interconnect_0_hex1_s1_readdata,                        --                                                     .readdata
			hex1_s1_writedata                                          => mm_interconnect_0_hex1_s1_writedata,                       --                                                     .writedata
			hex1_s1_chipselect                                         => mm_interconnect_0_hex1_s1_chipselect,                      --                                                     .chipselect
			hex2_s1_address                                            => mm_interconnect_0_hex2_s1_address,                         --                                              hex2_s1.address
			hex2_s1_write                                              => mm_interconnect_0_hex2_s1_write,                           --                                                     .write
			hex2_s1_readdata                                           => mm_interconnect_0_hex2_s1_readdata,                        --                                                     .readdata
			hex2_s1_writedata                                          => mm_interconnect_0_hex2_s1_writedata,                       --                                                     .writedata
			hex2_s1_chipselect                                         => mm_interconnect_0_hex2_s1_chipselect,                      --                                                     .chipselect
			hex3_s1_address                                            => mm_interconnect_0_hex3_s1_address,                         --                                              hex3_s1.address
			hex3_s1_write                                              => mm_interconnect_0_hex3_s1_write,                           --                                                     .write
			hex3_s1_readdata                                           => mm_interconnect_0_hex3_s1_readdata,                        --                                                     .readdata
			hex3_s1_writedata                                          => mm_interconnect_0_hex3_s1_writedata,                       --                                                     .writedata
			hex3_s1_chipselect                                         => mm_interconnect_0_hex3_s1_chipselect,                      --                                                     .chipselect
			hex4_s1_address                                            => mm_interconnect_0_hex4_s1_address,                         --                                              hex4_s1.address
			hex4_s1_write                                              => mm_interconnect_0_hex4_s1_write,                           --                                                     .write
			hex4_s1_readdata                                           => mm_interconnect_0_hex4_s1_readdata,                        --                                                     .readdata
			hex4_s1_writedata                                          => mm_interconnect_0_hex4_s1_writedata,                       --                                                     .writedata
			hex4_s1_chipselect                                         => mm_interconnect_0_hex4_s1_chipselect,                      --                                                     .chipselect
			hex5_s1_address                                            => mm_interconnect_0_hex5_s1_address,                         --                                              hex5_s1.address
			hex5_s1_write                                              => mm_interconnect_0_hex5_s1_write,                           --                                                     .write
			hex5_s1_readdata                                           => mm_interconnect_0_hex5_s1_readdata,                        --                                                     .readdata
			hex5_s1_writedata                                          => mm_interconnect_0_hex5_s1_writedata,                       --                                                     .writedata
			hex5_s1_chipselect                                         => mm_interconnect_0_hex5_s1_chipselect,                      --                                                     .chipselect
			jtag_uart_avalon_jtag_slave_address                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                          jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                     .write
			jtag_uart_avalon_jtag_slave_read                           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                     .read
			jtag_uart_avalon_jtag_slave_readdata                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                     .readdata
			jtag_uart_avalon_jtag_slave_writedata                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                     .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                     .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                     .chipselect
			led_s1_address                                             => mm_interconnect_0_led_s1_address,                          --                                               led_s1.address
			led_s1_write                                               => mm_interconnect_0_led_s1_write,                            --                                                     .write
			led_s1_readdata                                            => mm_interconnect_0_led_s1_readdata,                         --                                                     .readdata
			led_s1_writedata                                           => mm_interconnect_0_led_s1_writedata,                        --                                                     .writedata
			led_s1_chipselect                                          => mm_interconnect_0_led_s1_chipselect,                       --                                                     .chipselect
			onchip_memory_s1_address                                   => mm_interconnect_0_onchip_memory_s1_address,                --                                     onchip_memory_s1.address
			onchip_memory_s1_write                                     => mm_interconnect_0_onchip_memory_s1_write,                  --                                                     .write
			onchip_memory_s1_readdata                                  => mm_interconnect_0_onchip_memory_s1_readdata,               --                                                     .readdata
			onchip_memory_s1_writedata                                 => mm_interconnect_0_onchip_memory_s1_writedata,              --                                                     .writedata
			onchip_memory_s1_byteenable                                => mm_interconnect_0_onchip_memory_s1_byteenable,             --                                                     .byteenable
			onchip_memory_s1_chipselect                                => mm_interconnect_0_onchip_memory_s1_chipselect,             --                                                     .chipselect
			onchip_memory_s1_clken                                     => mm_interconnect_0_onchip_memory_s1_clken,                  --                                                     .clken
			sdram_s1_address                                           => mm_interconnect_0_sdram_s1_address,                        --                                             sdram_s1.address
			sdram_s1_write                                             => mm_interconnect_0_sdram_s1_write,                          --                                                     .write
			sdram_s1_read                                              => mm_interconnect_0_sdram_s1_read,                           --                                                     .read
			sdram_s1_readdata                                          => mm_interconnect_0_sdram_s1_readdata,                       --                                                     .readdata
			sdram_s1_writedata                                         => mm_interconnect_0_sdram_s1_writedata,                      --                                                     .writedata
			sdram_s1_byteenable                                        => mm_interconnect_0_sdram_s1_byteenable,                     --                                                     .byteenable
			sdram_s1_readdatavalid                                     => mm_interconnect_0_sdram_s1_readdatavalid,                  --                                                     .readdatavalid
			sdram_s1_waitrequest                                       => mm_interconnect_0_sdram_s1_waitrequest,                    --                                                     .waitrequest
			sdram_s1_chipselect                                        => mm_interconnect_0_sdram_s1_chipselect,                     --                                                     .chipselect
			switch_s1_address                                          => mm_interconnect_0_switch_s1_address,                       --                                            switch_s1.address
			switch_s1_readdata                                         => mm_interconnect_0_switch_s1_readdata,                      --                                                     .readdata
			sys_timer_s1_address                                       => mm_interconnect_0_sys_timer_s1_address,                    --                                         sys_timer_s1.address
			sys_timer_s1_write                                         => mm_interconnect_0_sys_timer_s1_write,                      --                                                     .write
			sys_timer_s1_readdata                                      => mm_interconnect_0_sys_timer_s1_readdata,                   --                                                     .readdata
			sys_timer_s1_writedata                                     => mm_interconnect_0_sys_timer_s1_writedata,                  --                                                     .writedata
			sys_timer_s1_chipselect                                    => mm_interconnect_0_sys_timer_s1_chipselect                  --                                                     .chipselect
		);

	irq_mapper : component platform_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                    --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	rst_controller : component platform_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component platform_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_debug_reset_request_reset,      -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component platform_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sys_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_timer_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_hex0_s1_write_ports_inv <= not mm_interconnect_0_hex0_s1_write;

	mm_interconnect_0_hex1_s1_write_ports_inv <= not mm_interconnect_0_hex1_s1_write;

	mm_interconnect_0_hex2_s1_write_ports_inv <= not mm_interconnect_0_hex2_s1_write;

	mm_interconnect_0_hex3_s1_write_ports_inv <= not mm_interconnect_0_hex3_s1_write;

	mm_interconnect_0_hex4_s1_write_ports_inv <= not mm_interconnect_0_hex4_s1_write;

	mm_interconnect_0_hex5_s1_write_ports_inv <= not mm_interconnect_0_hex5_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of platform
