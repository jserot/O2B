-- nios_128k_extended.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_128k_extended is
	port (
		button_external_connection_export : in  std_logic_vector(1 downto 0) := (others => '0'); -- button_external_connection.export
		clk_clk                           : in  std_logic                    := '0';             --                        clk.clk
		hex0_external_connection_export   : out std_logic_vector(7 downto 0);                    --   hex0_external_connection.export
		hex1_external_connection_export   : out std_logic_vector(7 downto 0);                    --   hex1_external_connection.export
		hex2_external_connection_export   : out std_logic_vector(7 downto 0);                    --   hex2_external_connection.export
		hex3_external_connection_export   : out std_logic_vector(7 downto 0);                    --   hex3_external_connection.export
		hex4_external_connection_export   : out std_logic_vector(7 downto 0);                    --   hex4_external_connection.export
		hex5_external_connection_export   : out std_logic_vector(7 downto 0);                    --   hex5_external_connection.export
		led_external_connection_export    : out std_logic_vector(9 downto 0);                    --    led_external_connection.export
		reset_reset_n                     : in  std_logic                    := '0';             --                      reset.reset_n
		switch_external_connection_export : in  std_logic_vector(9 downto 0) := (others => '0')  -- switch_external_connection.export
	);
end entity nios_128k_extended;

architecture rtl of nios_128k_extended is
	component nios_128k_extended_button is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component nios_128k_extended_button;

	component nios_128k_extended_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(18 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_multi_done                     : in  std_logic                     := 'X';             -- done
			E_ci_multi_clk_en                   : out std_logic;                                        -- clk_en
			E_ci_multi_start                    : out std_logic;                                        -- start
			E_ci_result                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                              : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                              : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                              : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                              : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                         : out std_logic;                                        -- readra
			D_ci_readrb                         : out std_logic;                                        -- readrb
			D_ci_writerc                        : out std_logic;                                        -- writerc
			E_ci_dataa                          : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                          : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                    : out std_logic;                                        -- clk
			E_ci_multi_reset                    : out std_logic;                                        -- reset
			E_ci_multi_reset_req                : out std_logic;                                        -- reset_req
			W_ci_estatus                        : out std_logic;                                        -- estatus
			W_ci_ipending                       : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component nios_128k_extended_cpu;

	component avs_gcd is
		port (
			avs_s0_address   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avs_s0_read      : in  std_logic                     := 'X';             -- read
			avs_s0_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write     : in  std_logic                     := 'X';             -- write
			avs_s0_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_clk        : in  std_logic                     := 'X';             -- clk
			reset_reset      : in  std_logic                     := 'X'              -- reset
		);
	end component avs_gcd;

	component custom_gcd is
		port (
			clk_en : in  std_logic                     := 'X';             -- clk_en
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			result : out std_logic_vector(31 downto 0);                    -- result
			clk    : in  std_logic                     := 'X';             -- clk
			reset  : in  std_logic                     := 'X'              -- reset
		);
	end component custom_gcd;

	component nios_128k_extended_hex0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios_128k_extended_hex0;

	component nios_128k_extended_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_128k_extended_jtag_uart;

	component nios_128k_extended_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component nios_128k_extended_led;

	component nios_128k_extended_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios_128k_extended_onchip_memory;

	component nios_128k_extended_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component nios_128k_extended_switch;

	component nios_128k_extended_sys_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_128k_extended_sys_id;

	component nios_128k_extended_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_128k_extended_timer;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X')  -- multi_c
		);
	end component altera_customins_master_translator;

	component nios_128k_extended_cpu_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result      : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra      : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb      : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc     : in  std_logic                     := 'X';             -- writerc
			ci_slave_a           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus     : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk         : in  std_logic                     := 'X';             -- clk
			ci_slave_reset       : in  std_logic                     := 'X';             -- reset
			ci_slave_clken       : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req   : in  std_logic                     := 'X';             -- reset_req
			ci_slave_start       : in  std_logic                     := 'X';             -- start
			ci_slave_done        : out std_logic;                                        -- done
			ci_master0_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra    : out std_logic;                                        -- readra
			ci_master0_readrb    : out std_logic;                                        -- readrb
			ci_master0_writerc   : out std_logic;                                        -- writerc
			ci_master0_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus   : out std_logic;                                        -- estatus
			ci_master0_clk       : out std_logic;                                        -- clk
			ci_master0_reset     : out std_logic;                                        -- reset
			ci_master0_clken     : out std_logic;                                        -- clk_en
			ci_master0_reset_req : out std_logic;                                        -- reset_req
			ci_master0_start     : out std_logic;                                        -- start
			ci_master0_done      : in  std_logic                     := 'X'              -- done
		);
	end component nios_128k_extended_cpu_custom_instruction_master_multi_xconnect;

	component altera_customins_slave_translator is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic;                                        -- done
			ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_clk       : out std_logic;                                        -- clk
			ci_master_clken     : out std_logic;                                        -- clk_en
			ci_master_reset     : out std_logic;                                        -- reset
			ci_master_start     : out std_logic;                                        -- start
			ci_master_done      : in  std_logic                     := 'X';             -- done
			ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master_readra    : out std_logic;                                        -- readra
			ci_master_readrb    : out std_logic;                                        -- readrb
			ci_master_writerc   : out std_logic;                                        -- writerc
			ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus   : out std_logic;                                        -- estatus
			ci_master_reset_req : out std_logic                                         -- reset_req
		);
	end component altera_customins_slave_translator;

	component nios_128k_extended_mm_interconnect_0 is
		port (
			clk_clk_clk                             : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                 : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address          : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			button_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			button_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			gcd_cc_s0_address                       : out std_logic_vector(3 downto 0);                     -- address
			gcd_cc_s0_write                         : out std_logic;                                        -- write
			gcd_cc_s0_read                          : out std_logic;                                        -- read
			gcd_cc_s0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			gcd_cc_s0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			hex0_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			hex0_s1_write                           : out std_logic;                                        -- write
			hex0_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex0_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex0_s1_chipselect                      : out std_logic;                                        -- chipselect
			hex1_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			hex1_s1_write                           : out std_logic;                                        -- write
			hex1_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex1_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex1_s1_chipselect                      : out std_logic;                                        -- chipselect
			hex2_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			hex2_s1_write                           : out std_logic;                                        -- write
			hex2_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex2_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex2_s1_chipselect                      : out std_logic;                                        -- chipselect
			hex3_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			hex3_s1_write                           : out std_logic;                                        -- write
			hex3_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex3_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex3_s1_chipselect                      : out std_logic;                                        -- chipselect
			hex4_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			hex4_s1_write                           : out std_logic;                                        -- write
			hex4_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex4_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex4_s1_chipselect                      : out std_logic;                                        -- chipselect
			hex5_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			hex5_s1_write                           : out std_logic;                                        -- write
			hex5_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex5_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex5_s1_chipselect                      : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			led_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                            : out std_logic;                                        -- write
			led_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                       : out std_logic;                                        -- chipselect
			onchip_memory_s1_address                : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory_s1_write                  : out std_logic;                                        -- write
			onchip_memory_s1_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect             : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                  : out std_logic;                                        -- clken
			switch_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_id_control_slave_address            : out std_logic_vector(0 downto 0);                     -- address
			sys_id_control_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                        : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                          : out std_logic;                                        -- write
			timer_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                     : out std_logic                                         -- chipselect
		);
	end component nios_128k_extended_mm_interconnect_0;

	component nios_128k_extended_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_128k_extended_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_custom_instruction_master_readra                                   : std_logic;                     -- cpu:D_ci_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	signal cpu_custom_instruction_master_a                                        : std_logic_vector(4 downto 0);  -- cpu:D_ci_a -> cpu_custom_instruction_master_translator:ci_slave_a
	signal cpu_custom_instruction_master_b                                        : std_logic_vector(4 downto 0);  -- cpu:D_ci_b -> cpu_custom_instruction_master_translator:ci_slave_b
	signal cpu_custom_instruction_master_c                                        : std_logic_vector(4 downto 0);  -- cpu:D_ci_c -> cpu_custom_instruction_master_translator:ci_slave_c
	signal cpu_custom_instruction_master_readrb                                   : std_logic;                     -- cpu:D_ci_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	signal cpu_custom_instruction_master_clk                                      : std_logic;                     -- cpu:E_ci_multi_clock -> cpu_custom_instruction_master_translator:ci_slave_multi_clk
	signal cpu_custom_instruction_master_ipending                                 : std_logic_vector(31 downto 0); -- cpu:W_ci_ipending -> cpu_custom_instruction_master_translator:ci_slave_ipending
	signal cpu_custom_instruction_master_start                                    : std_logic;                     -- cpu:E_ci_multi_start -> cpu_custom_instruction_master_translator:ci_slave_multi_start
	signal cpu_custom_instruction_master_reset_req                                : std_logic;                     -- cpu:E_ci_multi_reset_req -> cpu_custom_instruction_master_translator:ci_slave_multi_reset_req
	signal cpu_custom_instruction_master_done                                     : std_logic;                     -- cpu_custom_instruction_master_translator:ci_slave_multi_done -> cpu:E_ci_multi_done
	signal cpu_custom_instruction_master_n                                        : std_logic_vector(7 downto 0);  -- cpu:D_ci_n -> cpu_custom_instruction_master_translator:ci_slave_n
	signal cpu_custom_instruction_master_result                                   : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_result
	signal cpu_custom_instruction_master_estatus                                  : std_logic;                     -- cpu:W_ci_estatus -> cpu_custom_instruction_master_translator:ci_slave_estatus
	signal cpu_custom_instruction_master_clk_en                                   : std_logic;                     -- cpu:E_ci_multi_clk_en -> cpu_custom_instruction_master_translator:ci_slave_multi_clken
	signal cpu_custom_instruction_master_datab                                    : std_logic_vector(31 downto 0); -- cpu:E_ci_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	signal cpu_custom_instruction_master_dataa                                    : std_logic_vector(31 downto 0); -- cpu:E_ci_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	signal cpu_custom_instruction_master_reset                                    : std_logic;                     -- cpu:E_ci_multi_reset -> cpu_custom_instruction_master_translator:ci_slave_multi_reset
	signal cpu_custom_instruction_master_writerc                                  : std_logic;                     -- cpu:D_ci_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	signal cpu_custom_instruction_master_translator_multi_ci_master_readra        : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_readra -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal cpu_custom_instruction_master_translator_multi_ci_master_a             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_a -> cpu_custom_instruction_master_multi_xconnect:ci_slave_a
	signal cpu_custom_instruction_master_translator_multi_ci_master_b             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_b -> cpu_custom_instruction_master_multi_xconnect:ci_slave_b
	signal cpu_custom_instruction_master_translator_multi_ci_master_clk           : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_clk -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal cpu_custom_instruction_master_translator_multi_ci_master_readrb        : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal cpu_custom_instruction_master_translator_multi_ci_master_c             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_c -> cpu_custom_instruction_master_multi_xconnect:ci_slave_c
	signal cpu_custom_instruction_master_translator_multi_ci_master_start         : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_start -> cpu_custom_instruction_master_multi_xconnect:ci_slave_start
	signal cpu_custom_instruction_master_translator_multi_ci_master_reset_req     : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	signal cpu_custom_instruction_master_translator_multi_ci_master_done          : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_custom_instruction_master_translator:multi_ci_master_done
	signal cpu_custom_instruction_master_translator_multi_ci_master_n             : std_logic_vector(7 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_n -> cpu_custom_instruction_master_multi_xconnect:ci_slave_n
	signal cpu_custom_instruction_master_translator_multi_ci_master_result        : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:multi_ci_master_result
	signal cpu_custom_instruction_master_translator_multi_ci_master_clk_en        : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_clken -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal cpu_custom_instruction_master_translator_multi_ci_master_datab         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:multi_ci_master_datab -> cpu_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal cpu_custom_instruction_master_translator_multi_ci_master_dataa         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal cpu_custom_instruction_master_translator_multi_ci_master_reset         : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_reset -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal cpu_custom_instruction_master_translator_multi_ci_master_writerc       : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_readra         : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb         : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_clk            : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_start          : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req      : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_done           : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_custom_instruction_master_multi_xconnect:ci_master0_done
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_multi_xconnect:ci_master0_result
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus        : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en         : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_reset          : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc        : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- gcd_ci:result -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk    : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_clk -> gcd_ci:clk
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_clken -> gcd_ci:clk_en
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab  : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_datab -> gcd_ci:datab
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> gcd_ci:dataa
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_start  : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_start -> gcd_ci:start
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset  : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset -> gcd_ci:reset
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_done   : std_logic;                     -- gcd_ci:done -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal cpu_data_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                            : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                : std_logic_vector(18 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                             : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                   : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                  : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                              : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                         : std_logic_vector(18 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                            : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect               : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                 : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest              : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                     : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                    : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sys_id_control_slave_readdata                        : std_logic_vector(31 downto 0); -- sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	signal mm_interconnect_0_sys_id_control_slave_address                         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                         : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                      : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                      : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                             : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                            : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_gcd_cc_s0_readdata                                   : std_logic_vector(31 downto 0); -- gcd_cc:avs_s0_readdata -> mm_interconnect_0:gcd_cc_s0_readdata
	signal mm_interconnect_0_gcd_cc_s0_address                                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:gcd_cc_s0_address -> gcd_cc:avs_s0_address
	signal mm_interconnect_0_gcd_cc_s0_read                                       : std_logic;                     -- mm_interconnect_0:gcd_cc_s0_read -> gcd_cc:avs_s0_read
	signal mm_interconnect_0_gcd_cc_s0_write                                      : std_logic;                     -- mm_interconnect_0:gcd_cc_s0_write -> gcd_cc:avs_s0_write
	signal mm_interconnect_0_gcd_cc_s0_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:gcd_cc_s0_writedata -> gcd_cc:avs_s0_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                            : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                             : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                               : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                               : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_button_s1_readdata                                   : std_logic_vector(31 downto 0); -- button:readdata -> mm_interconnect_0:button_s1_readdata
	signal mm_interconnect_0_button_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_s1_address -> button:address
	signal mm_interconnect_0_switch_s1_readdata                                   : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_led_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                                      : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                                         : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_hex0_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	signal mm_interconnect_0_hex0_s1_readdata                                     : std_logic_vector(31 downto 0); -- hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	signal mm_interconnect_0_hex0_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex0_s1_address -> hex0:address
	signal mm_interconnect_0_hex0_s1_write                                        : std_logic;                     -- mm_interconnect_0:hex0_s1_write -> mm_interconnect_0_hex0_s1_write:in
	signal mm_interconnect_0_hex0_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	signal mm_interconnect_0_hex1_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	signal mm_interconnect_0_hex1_s1_readdata                                     : std_logic_vector(31 downto 0); -- hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	signal mm_interconnect_0_hex1_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex1_s1_address -> hex1:address
	signal mm_interconnect_0_hex1_s1_write                                        : std_logic;                     -- mm_interconnect_0:hex1_s1_write -> mm_interconnect_0_hex1_s1_write:in
	signal mm_interconnect_0_hex1_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	signal mm_interconnect_0_hex2_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	signal mm_interconnect_0_hex2_s1_readdata                                     : std_logic_vector(31 downto 0); -- hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	signal mm_interconnect_0_hex2_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex2_s1_address -> hex2:address
	signal mm_interconnect_0_hex2_s1_write                                        : std_logic;                     -- mm_interconnect_0:hex2_s1_write -> mm_interconnect_0_hex2_s1_write:in
	signal mm_interconnect_0_hex2_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	signal mm_interconnect_0_hex3_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	signal mm_interconnect_0_hex3_s1_readdata                                     : std_logic_vector(31 downto 0); -- hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	signal mm_interconnect_0_hex3_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex3_s1_address -> hex3:address
	signal mm_interconnect_0_hex3_s1_write                                        : std_logic;                     -- mm_interconnect_0:hex3_s1_write -> mm_interconnect_0_hex3_s1_write:in
	signal mm_interconnect_0_hex3_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	signal mm_interconnect_0_hex4_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	signal mm_interconnect_0_hex4_s1_readdata                                     : std_logic_vector(31 downto 0); -- hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	signal mm_interconnect_0_hex4_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex4_s1_address -> hex4:address
	signal mm_interconnect_0_hex4_s1_write                                        : std_logic;                     -- mm_interconnect_0:hex4_s1_write -> mm_interconnect_0_hex4_s1_write:in
	signal mm_interconnect_0_hex4_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	signal mm_interconnect_0_hex5_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	signal mm_interconnect_0_hex5_s1_readdata                                     : std_logic_vector(31 downto 0); -- hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	signal mm_interconnect_0_hex5_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex5_s1_address -> hex5:address
	signal mm_interconnect_0_hex5_s1_write                                        : std_logic;                     -- mm_interconnect_0:hex5_s1_write -> mm_interconnect_0_hex5_s1_write:in
	signal mm_interconnect_0_hex5_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	signal mm_interconnect_0_timer_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                                    : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_0:timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                                     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_s1_address -> timer:address
	signal mm_interconnect_0_timer_s1_write                                       : std_logic;                     -- mm_interconnect_0:timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_s1_writedata -> timer:writedata
	signal irq_mapper_receiver0_irq                                               : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                               : std_logic;                     -- timer:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                         : std_logic;                     -- rst_controller:reset_out -> [gcd_cc:reset_reset, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                     : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                                : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv           : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_hex0_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_hex0_s1_write:inv -> hex0:write_n
	signal mm_interconnect_0_hex1_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_hex1_s1_write:inv -> hex1:write_n
	signal mm_interconnect_0_hex2_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_hex2_s1_write:inv -> hex2:write_n
	signal mm_interconnect_0_hex3_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_hex3_s1_write:inv -> hex3:write_n
	signal mm_interconnect_0_hex4_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_hex4_s1_write:inv -> hex4:write_n
	signal mm_interconnect_0_hex5_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_hex5_s1_write:inv -> hex5:write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [button:reset_n, cpu:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, jtag_uart:rst_n, led:reset_n, switch:reset_n, sys_id:reset_n, timer:reset_n]

begin

	button : component nios_128k_extended_button
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_button_s1_readdata,     --                    .readdata
			in_port  => button_external_connection_export         -- external_connection.export
		);

	cpu : component nios_128k_extended_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			E_ci_multi_done                     => cpu_custom_instruction_master_done,                -- custom_instruction_master.done
			E_ci_multi_clk_en                   => cpu_custom_instruction_master_clk_en,              --                          .clk_en
			E_ci_multi_start                    => cpu_custom_instruction_master_start,               --                          .start
			E_ci_result                         => cpu_custom_instruction_master_result,              --                          .result
			D_ci_a                              => cpu_custom_instruction_master_a,                   --                          .a
			D_ci_b                              => cpu_custom_instruction_master_b,                   --                          .b
			D_ci_c                              => cpu_custom_instruction_master_c,                   --                          .c
			D_ci_n                              => cpu_custom_instruction_master_n,                   --                          .n
			D_ci_readra                         => cpu_custom_instruction_master_readra,              --                          .readra
			D_ci_readrb                         => cpu_custom_instruction_master_readrb,              --                          .readrb
			D_ci_writerc                        => cpu_custom_instruction_master_writerc,             --                          .writerc
			E_ci_dataa                          => cpu_custom_instruction_master_dataa,               --                          .dataa
			E_ci_datab                          => cpu_custom_instruction_master_datab,               --                          .datab
			E_ci_multi_clock                    => cpu_custom_instruction_master_clk,                 --                          .clk
			E_ci_multi_reset                    => cpu_custom_instruction_master_reset,               --                          .reset
			E_ci_multi_reset_req                => cpu_custom_instruction_master_reset_req,           --                          .reset_req
			W_ci_estatus                        => cpu_custom_instruction_master_estatus,             --                          .estatus
			W_ci_ipending                       => cpu_custom_instruction_master_ipending             --                          .ipending
		);

	gcd_cc : component avs_gcd
		port map (
			avs_s0_address   => mm_interconnect_0_gcd_cc_s0_address,   --    s0.address
			avs_s0_read      => mm_interconnect_0_gcd_cc_s0_read,      --      .read
			avs_s0_readdata  => mm_interconnect_0_gcd_cc_s0_readdata,  --      .readdata
			avs_s0_write     => mm_interconnect_0_gcd_cc_s0_write,     --      .write
			avs_s0_writedata => mm_interconnect_0_gcd_cc_s0_writedata, --      .writedata
			clock_clk        => clk_clk,                               -- clock.clk
			reset_reset      => rst_controller_reset_out_reset         -- reset.reset
		);

	gcd_ci : component custom_gcd
		port map (
			clk_en => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, -- nios_custom_instruction_slave.clk_en
			start  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_start,  --                              .start
			done   => cpu_custom_instruction_master_multi_slave_translator0_ci_master_done,   --                              .done
			dataa  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --                              .dataa
			datab  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --                              .datab
			result => cpu_custom_instruction_master_multi_slave_translator0_ci_master_result, --                              .result
			clk    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --                              .clk
			reset  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset   --                              .reset
		);

	hex0 : component nios_128k_extended_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex0_s1_readdata,        --                    .readdata
			out_port   => hex0_external_connection_export            -- external_connection.export
		);

	hex1 : component nios_128k_extended_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex1_s1_readdata,        --                    .readdata
			out_port   => hex1_external_connection_export            -- external_connection.export
		);

	hex2 : component nios_128k_extended_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex2_s1_readdata,        --                    .readdata
			out_port   => hex2_external_connection_export            -- external_connection.export
		);

	hex3 : component nios_128k_extended_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex3_s1_readdata,        --                    .readdata
			out_port   => hex3_external_connection_export            -- external_connection.export
		);

	hex4 : component nios_128k_extended_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex4_s1_readdata,        --                    .readdata
			out_port   => hex4_external_connection_export            -- external_connection.export
		);

	hex5 : component nios_128k_extended_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex5_s1_readdata,        --                    .readdata
			out_port   => hex5_external_connection_export            -- external_connection.export
		);

	jtag_uart : component nios_128k_extended_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	led : component nios_128k_extended_led
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	onchip_memory : component nios_128k_extended_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req             --       .reset_req
		);

	switch : component nios_128k_extended_switch
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_external_connection_export         -- external_connection.export
		);

	sys_id : component nios_128k_extended_sys_id
		port map (
			clock    => clk_clk,                                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_sys_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sys_id_control_slave_address(0)  --              .address
		);

	timer : component nios_128k_extended_timer
		port map (
			clk        => clk_clk,                                    --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                    --   irq.irq
		);

	cpu_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa            => cpu_custom_instruction_master_dataa,                                --        ci_slave.dataa
			ci_slave_datab            => cpu_custom_instruction_master_datab,                                --                .datab
			ci_slave_result           => cpu_custom_instruction_master_result,                               --                .result
			ci_slave_n                => cpu_custom_instruction_master_n,                                    --                .n
			ci_slave_readra           => cpu_custom_instruction_master_readra,                               --                .readra
			ci_slave_readrb           => cpu_custom_instruction_master_readrb,                               --                .readrb
			ci_slave_writerc          => cpu_custom_instruction_master_writerc,                              --                .writerc
			ci_slave_a                => cpu_custom_instruction_master_a,                                    --                .a
			ci_slave_b                => cpu_custom_instruction_master_b,                                    --                .b
			ci_slave_c                => cpu_custom_instruction_master_c,                                    --                .c
			ci_slave_ipending         => cpu_custom_instruction_master_ipending,                             --                .ipending
			ci_slave_estatus          => cpu_custom_instruction_master_estatus,                              --                .estatus
			ci_slave_multi_clk        => cpu_custom_instruction_master_clk,                                  --                .clk
			ci_slave_multi_reset      => cpu_custom_instruction_master_reset,                                --                .reset
			ci_slave_multi_clken      => cpu_custom_instruction_master_clk_en,                               --                .clk_en
			ci_slave_multi_reset_req  => cpu_custom_instruction_master_reset_req,                            --                .reset_req
			ci_slave_multi_start      => cpu_custom_instruction_master_start,                                --                .start
			ci_slave_multi_done       => cpu_custom_instruction_master_done,                                 --                .done
			comb_ci_master_dataa      => open,                                                               --  comb_ci_master.dataa
			comb_ci_master_datab      => open,                                                               --                .datab
			comb_ci_master_result     => open,                                                               --                .result
			comb_ci_master_n          => open,                                                               --                .n
			comb_ci_master_readra     => open,                                                               --                .readra
			comb_ci_master_readrb     => open,                                                               --                .readrb
			comb_ci_master_writerc    => open,                                                               --                .writerc
			comb_ci_master_a          => open,                                                               --                .a
			comb_ci_master_b          => open,                                                               --                .b
			comb_ci_master_c          => open,                                                               --                .c
			comb_ci_master_ipending   => open,                                                               --                .ipending
			comb_ci_master_estatus    => open,                                                               --                .estatus
			multi_ci_master_clk       => cpu_custom_instruction_master_translator_multi_ci_master_clk,       -- multi_ci_master.clk
			multi_ci_master_reset     => cpu_custom_instruction_master_translator_multi_ci_master_reset,     --                .reset
			multi_ci_master_clken     => cpu_custom_instruction_master_translator_multi_ci_master_clk_en,    --                .clk_en
			multi_ci_master_reset_req => cpu_custom_instruction_master_translator_multi_ci_master_reset_req, --                .reset_req
			multi_ci_master_start     => cpu_custom_instruction_master_translator_multi_ci_master_start,     --                .start
			multi_ci_master_done      => cpu_custom_instruction_master_translator_multi_ci_master_done,      --                .done
			multi_ci_master_dataa     => cpu_custom_instruction_master_translator_multi_ci_master_dataa,     --                .dataa
			multi_ci_master_datab     => cpu_custom_instruction_master_translator_multi_ci_master_datab,     --                .datab
			multi_ci_master_result    => cpu_custom_instruction_master_translator_multi_ci_master_result,    --                .result
			multi_ci_master_n         => cpu_custom_instruction_master_translator_multi_ci_master_n,         --                .n
			multi_ci_master_readra    => cpu_custom_instruction_master_translator_multi_ci_master_readra,    --                .readra
			multi_ci_master_readrb    => cpu_custom_instruction_master_translator_multi_ci_master_readrb,    --                .readrb
			multi_ci_master_writerc   => cpu_custom_instruction_master_translator_multi_ci_master_writerc,   --                .writerc
			multi_ci_master_a         => cpu_custom_instruction_master_translator_multi_ci_master_a,         --                .a
			multi_ci_master_b         => cpu_custom_instruction_master_translator_multi_ci_master_b,         --                .b
			multi_ci_master_c         => cpu_custom_instruction_master_translator_multi_ci_master_c,         --                .c
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                                 --     (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                                 --     (terminated)
			ci_slave_multi_result     => open,                                                               --     (terminated)
			ci_slave_multi_n          => "00000000",                                                         --     (terminated)
			ci_slave_multi_readra     => '0',                                                                --     (terminated)
			ci_slave_multi_readrb     => '0',                                                                --     (terminated)
			ci_slave_multi_writerc    => '0',                                                                --     (terminated)
			ci_slave_multi_a          => "00000",                                                            --     (terminated)
			ci_slave_multi_b          => "00000",                                                            --     (terminated)
			ci_slave_multi_c          => "00000"                                                             --     (terminated)
		);

	cpu_custom_instruction_master_multi_xconnect : component nios_128k_extended_cpu_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa       => cpu_custom_instruction_master_translator_multi_ci_master_dataa,     --   ci_slave.dataa
			ci_slave_datab       => cpu_custom_instruction_master_translator_multi_ci_master_datab,     --           .datab
			ci_slave_result      => cpu_custom_instruction_master_translator_multi_ci_master_result,    --           .result
			ci_slave_n           => cpu_custom_instruction_master_translator_multi_ci_master_n,         --           .n
			ci_slave_readra      => cpu_custom_instruction_master_translator_multi_ci_master_readra,    --           .readra
			ci_slave_readrb      => cpu_custom_instruction_master_translator_multi_ci_master_readrb,    --           .readrb
			ci_slave_writerc     => cpu_custom_instruction_master_translator_multi_ci_master_writerc,   --           .writerc
			ci_slave_a           => cpu_custom_instruction_master_translator_multi_ci_master_a,         --           .a
			ci_slave_b           => cpu_custom_instruction_master_translator_multi_ci_master_b,         --           .b
			ci_slave_c           => cpu_custom_instruction_master_translator_multi_ci_master_c,         --           .c
			ci_slave_ipending    => open,                                                               --           .ipending
			ci_slave_estatus     => open,                                                               --           .estatus
			ci_slave_clk         => cpu_custom_instruction_master_translator_multi_ci_master_clk,       --           .clk
			ci_slave_reset       => cpu_custom_instruction_master_translator_multi_ci_master_reset,     --           .reset
			ci_slave_clken       => cpu_custom_instruction_master_translator_multi_ci_master_clk_en,    --           .clk_en
			ci_slave_reset_req   => cpu_custom_instruction_master_translator_multi_ci_master_reset_req, --           .reset_req
			ci_slave_start       => cpu_custom_instruction_master_translator_multi_ci_master_start,     --           .start
			ci_slave_done        => cpu_custom_instruction_master_translator_multi_ci_master_done,      --           .done
			ci_master0_dataa     => cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa,      -- ci_master0.dataa
			ci_master0_datab     => cpu_custom_instruction_master_multi_xconnect_ci_master0_datab,      --           .datab
			ci_master0_result    => cpu_custom_instruction_master_multi_xconnect_ci_master0_result,     --           .result
			ci_master0_n         => cpu_custom_instruction_master_multi_xconnect_ci_master0_n,          --           .n
			ci_master0_readra    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readra,     --           .readra
			ci_master0_readrb    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb,     --           .readrb
			ci_master0_writerc   => cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc,    --           .writerc
			ci_master0_a         => cpu_custom_instruction_master_multi_xconnect_ci_master0_a,          --           .a
			ci_master0_b         => cpu_custom_instruction_master_multi_xconnect_ci_master0_b,          --           .b
			ci_master0_c         => cpu_custom_instruction_master_multi_xconnect_ci_master0_c,          --           .c
			ci_master0_ipending  => cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending,   --           .ipending
			ci_master0_estatus   => cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus,    --           .estatus
			ci_master0_clk       => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk,        --           .clk
			ci_master0_reset     => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset,      --           .reset
			ci_master0_clken     => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en,     --           .clk_en
			ci_master0_reset_req => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req,  --           .reset_req
			ci_master0_start     => cpu_custom_instruction_master_multi_xconnect_ci_master0_start,      --           .start
			ci_master0_done      => cpu_custom_instruction_master_multi_xconnect_ci_master0_done        --           .done
		);

	cpu_custom_instruction_master_multi_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 8,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 0
		)
		port map (
			ci_slave_dataa      => cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => cpu_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => cpu_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => cpu_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => cpu_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => cpu_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => cpu_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => cpu_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk        => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken      => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset_req  => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req,      --          .reset_req
			ci_slave_reset      => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start      => cpu_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done       => cpu_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_clk       => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --          .clk_en
			ci_master_reset     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done      => cpu_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_n         => open,                                                                   -- (terminated)
			ci_master_readra    => open,                                                                   -- (terminated)
			ci_master_readrb    => open,                                                                   -- (terminated)
			ci_master_writerc   => open,                                                                   -- (terminated)
			ci_master_a         => open,                                                                   -- (terminated)
			ci_master_b         => open,                                                                   -- (terminated)
			ci_master_c         => open,                                                                   -- (terminated)
			ci_master_ipending  => open,                                                                   -- (terminated)
			ci_master_estatus   => open,                                                                   -- (terminated)
			ci_master_reset_req => open                                                                    -- (terminated)
		);

	mm_interconnect_0 : component nios_128k_extended_mm_interconnect_0
		port map (
			clk_clk_clk                             => clk_clk,                                                   --                         clk_clk.clk
			cpu_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                            -- cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                 => cpu_data_master_address,                                   --                 cpu_data_master.address
			cpu_data_master_waitrequest             => cpu_data_master_waitrequest,                               --                                .waitrequest
			cpu_data_master_byteenable              => cpu_data_master_byteenable,                                --                                .byteenable
			cpu_data_master_read                    => cpu_data_master_read,                                      --                                .read
			cpu_data_master_readdata                => cpu_data_master_readdata,                                  --                                .readdata
			cpu_data_master_write                   => cpu_data_master_write,                                     --                                .write
			cpu_data_master_writedata               => cpu_data_master_writedata,                                 --                                .writedata
			cpu_data_master_debugaccess             => cpu_data_master_debugaccess,                               --                                .debugaccess
			cpu_instruction_master_address          => cpu_instruction_master_address,                            --          cpu_instruction_master.address
			cpu_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                        --                                .waitrequest
			cpu_instruction_master_read             => cpu_instruction_master_read,                               --                                .read
			cpu_instruction_master_readdata         => cpu_instruction_master_readdata,                           --                                .readdata
			button_s1_address                       => mm_interconnect_0_button_s1_address,                       --                       button_s1.address
			button_s1_readdata                      => mm_interconnect_0_button_s1_readdata,                      --                                .readdata
			cpu_debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,             --             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                .write
			cpu_debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                .read
			cpu_debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                .readdata
			cpu_debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                .writedata
			cpu_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                .byteenable
			cpu_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                .waitrequest
			cpu_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                .debugaccess
			gcd_cc_s0_address                       => mm_interconnect_0_gcd_cc_s0_address,                       --                       gcd_cc_s0.address
			gcd_cc_s0_write                         => mm_interconnect_0_gcd_cc_s0_write,                         --                                .write
			gcd_cc_s0_read                          => mm_interconnect_0_gcd_cc_s0_read,                          --                                .read
			gcd_cc_s0_readdata                      => mm_interconnect_0_gcd_cc_s0_readdata,                      --                                .readdata
			gcd_cc_s0_writedata                     => mm_interconnect_0_gcd_cc_s0_writedata,                     --                                .writedata
			hex0_s1_address                         => mm_interconnect_0_hex0_s1_address,                         --                         hex0_s1.address
			hex0_s1_write                           => mm_interconnect_0_hex0_s1_write,                           --                                .write
			hex0_s1_readdata                        => mm_interconnect_0_hex0_s1_readdata,                        --                                .readdata
			hex0_s1_writedata                       => mm_interconnect_0_hex0_s1_writedata,                       --                                .writedata
			hex0_s1_chipselect                      => mm_interconnect_0_hex0_s1_chipselect,                      --                                .chipselect
			hex1_s1_address                         => mm_interconnect_0_hex1_s1_address,                         --                         hex1_s1.address
			hex1_s1_write                           => mm_interconnect_0_hex1_s1_write,                           --                                .write
			hex1_s1_readdata                        => mm_interconnect_0_hex1_s1_readdata,                        --                                .readdata
			hex1_s1_writedata                       => mm_interconnect_0_hex1_s1_writedata,                       --                                .writedata
			hex1_s1_chipselect                      => mm_interconnect_0_hex1_s1_chipselect,                      --                                .chipselect
			hex2_s1_address                         => mm_interconnect_0_hex2_s1_address,                         --                         hex2_s1.address
			hex2_s1_write                           => mm_interconnect_0_hex2_s1_write,                           --                                .write
			hex2_s1_readdata                        => mm_interconnect_0_hex2_s1_readdata,                        --                                .readdata
			hex2_s1_writedata                       => mm_interconnect_0_hex2_s1_writedata,                       --                                .writedata
			hex2_s1_chipselect                      => mm_interconnect_0_hex2_s1_chipselect,                      --                                .chipselect
			hex3_s1_address                         => mm_interconnect_0_hex3_s1_address,                         --                         hex3_s1.address
			hex3_s1_write                           => mm_interconnect_0_hex3_s1_write,                           --                                .write
			hex3_s1_readdata                        => mm_interconnect_0_hex3_s1_readdata,                        --                                .readdata
			hex3_s1_writedata                       => mm_interconnect_0_hex3_s1_writedata,                       --                                .writedata
			hex3_s1_chipselect                      => mm_interconnect_0_hex3_s1_chipselect,                      --                                .chipselect
			hex4_s1_address                         => mm_interconnect_0_hex4_s1_address,                         --                         hex4_s1.address
			hex4_s1_write                           => mm_interconnect_0_hex4_s1_write,                           --                                .write
			hex4_s1_readdata                        => mm_interconnect_0_hex4_s1_readdata,                        --                                .readdata
			hex4_s1_writedata                       => mm_interconnect_0_hex4_s1_writedata,                       --                                .writedata
			hex4_s1_chipselect                      => mm_interconnect_0_hex4_s1_chipselect,                      --                                .chipselect
			hex5_s1_address                         => mm_interconnect_0_hex5_s1_address,                         --                         hex5_s1.address
			hex5_s1_write                           => mm_interconnect_0_hex5_s1_write,                           --                                .write
			hex5_s1_readdata                        => mm_interconnect_0_hex5_s1_readdata,                        --                                .readdata
			hex5_s1_writedata                       => mm_interconnect_0_hex5_s1_writedata,                       --                                .writedata
			hex5_s1_chipselect                      => mm_interconnect_0_hex5_s1_chipselect,                      --                                .chipselect
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                .chipselect
			led_s1_address                          => mm_interconnect_0_led_s1_address,                          --                          led_s1.address
			led_s1_write                            => mm_interconnect_0_led_s1_write,                            --                                .write
			led_s1_readdata                         => mm_interconnect_0_led_s1_readdata,                         --                                .readdata
			led_s1_writedata                        => mm_interconnect_0_led_s1_writedata,                        --                                .writedata
			led_s1_chipselect                       => mm_interconnect_0_led_s1_chipselect,                       --                                .chipselect
			onchip_memory_s1_address                => mm_interconnect_0_onchip_memory_s1_address,                --                onchip_memory_s1.address
			onchip_memory_s1_write                  => mm_interconnect_0_onchip_memory_s1_write,                  --                                .write
			onchip_memory_s1_readdata               => mm_interconnect_0_onchip_memory_s1_readdata,               --                                .readdata
			onchip_memory_s1_writedata              => mm_interconnect_0_onchip_memory_s1_writedata,              --                                .writedata
			onchip_memory_s1_byteenable             => mm_interconnect_0_onchip_memory_s1_byteenable,             --                                .byteenable
			onchip_memory_s1_chipselect             => mm_interconnect_0_onchip_memory_s1_chipselect,             --                                .chipselect
			onchip_memory_s1_clken                  => mm_interconnect_0_onchip_memory_s1_clken,                  --                                .clken
			switch_s1_address                       => mm_interconnect_0_switch_s1_address,                       --                       switch_s1.address
			switch_s1_readdata                      => mm_interconnect_0_switch_s1_readdata,                      --                                .readdata
			sys_id_control_slave_address            => mm_interconnect_0_sys_id_control_slave_address,            --            sys_id_control_slave.address
			sys_id_control_slave_readdata           => mm_interconnect_0_sys_id_control_slave_readdata,           --                                .readdata
			timer_s1_address                        => mm_interconnect_0_timer_s1_address,                        --                        timer_s1.address
			timer_s1_write                          => mm_interconnect_0_timer_s1_write,                          --                                .write
			timer_s1_readdata                       => mm_interconnect_0_timer_s1_readdata,                       --                                .readdata
			timer_s1_writedata                      => mm_interconnect_0_timer_s1_writedata,                      --                                .writedata
			timer_s1_chipselect                     => mm_interconnect_0_timer_s1_chipselect                      --                                .chipselect
		);

	irq_mapper : component nios_128k_extended_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_hex0_s1_write_ports_inv <= not mm_interconnect_0_hex0_s1_write;

	mm_interconnect_0_hex1_s1_write_ports_inv <= not mm_interconnect_0_hex1_s1_write;

	mm_interconnect_0_hex2_s1_write_ports_inv <= not mm_interconnect_0_hex2_s1_write;

	mm_interconnect_0_hex3_s1_write_ports_inv <= not mm_interconnect_0_hex3_s1_write;

	mm_interconnect_0_hex4_s1_write_ports_inv <= not mm_interconnect_0_hex4_s1_write;

	mm_interconnect_0_hex5_s1_write_ports_inv <= not mm_interconnect_0_hex5_s1_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_128k_extended
